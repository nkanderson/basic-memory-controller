//////////////////////////////////////////////////////////////
// tc_mc_top.sv - Top level module for testing memory controller
//
// Author: Niklas Anderson (niklas2@pdx.edu)
// Date: Feb 26, 2025
//
// Description:
// ------------
// Top level module which instantiates the interface, memory
// controller, and the processor. Also generates the clock and
// reset signal in order to start the system.
//
////////////////////////////////////////////////////////////////

module tc_mc_top ();


endmodule
