//////////////////////////////////////////////////////////////
// processor.sv - Simulate a processor to test a memory controller
//
// Author: Niklas Anderson (niklas2@pdx.edu)
// Date: Feb 26, 2025
//
// Description:
// ------------
// Serves as a testbench for a memory controller module.
// Does this by simulating a processor.
//
////////////////////////////////////////////////////////////////

module processor();


endmodule
